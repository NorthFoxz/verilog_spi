module clock_sync()

endmodule